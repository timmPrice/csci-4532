module dfmult (
    input  wire a,
    input  wire b,
    input  wire addr,
    input  wire clk,
    output reg  q
);



endmodule




















