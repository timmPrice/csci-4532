module and(x, y, z)
    input x;
    input y;
    output z; 

    assign x&y=z;
endmodule
